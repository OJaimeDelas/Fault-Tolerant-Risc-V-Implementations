DEADC0B730001073
DEADC137EEF08093
DEADC1B7EEF10113
DEADC237EEF18193
DEADC2B7EEF20213
DEADC337EEF28293
DEADC3B7EEF30313
DEADC437EEF38393
DEADC4B7EEF40413
DEADC537EEF48493
DEADC5B7EEF50513
DEADC637EEF58593
DEADC6B7EEF60613
DEADC737EEF68693
DEADC7B7EEF70713
DEADC837EEF78793
DEADC8B7EEF80813
DEADC937EEF88893
DEADC9B7EEF90913
DEADCA37EEF98993
DEADCAB7EEFA0A13
DEADCB37EEFA8A93
DEADCBB7EEFB0B13
DEADCC37EEFB8B93
DEADCCB7EEFC0C13
DEADCD37EEFC8C93
DEADCDB7EEFD0D13
DEADCE37EEFD8D93
DEADCEB7EEFE0E13
DEADCF37EEFE8E93
DEADCFB7EEFF0F13
30401073EEFF8F93
3410107334001073
B000107334401073
B0301073B0201073
B0501073B0401073
B8001073B0601073
B8301073B8201073
B8501073B8401073
32301073B8601073
3250107332401073
7A00107332601073
5553031355555337
0000100F7C031073
0007866300000793
000000E700000097
000401370040006F
000011B700010113
F14027F34C818193
0000079300079C63
0000029302078263
0D00006F30529073
3052907322400293
00000793018000EF
22000293FE0792E3
0B00006F30529073
04B5506300100593
00058593000015B7
FFF5051340B10133
00001517FE051CE3
00052583B3450513
000007B7FE058EE3
0007886300078793
00000097F1402573
000007B7000000E7
0007866326878793
058080E700000097
FFDFF06F10500073
0000006F0000006F
00112823FE810113
00A1202300B12423
82E1AC2300100713
0007866300000793
000000E700000097
0005846300812583
010120837C60D073
0000806701810113
FF01011300008067
8501859300000613
0011262385018513
00000613640000EF
8501851300000593
850185137F0000EF
0E9000EF1C1000EF
84F1A42300100793
000005930FF0000F
54C000EF00000513
00000000171000EF
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0010031384C18293
00300E1300200393
01F0071300400E93
003006130062A023
0000001300000013
0000001300000013
0002AF0300000013
41CE8E3301EE8EB3
01C3F3B301D383B3
006393B300100693
406686B30AA3C393
00E3F3B3FE06DAE3
000000130072A023
0000001300000013
0000001300000013
0020039300100313
00400E9300300E13
F8061AE3FFF60613
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0100029300050F93
00060E6302567463
0005828300B60733
0055002300158593
FEE5E8E300150513
00008067000F8513
0035F39300357313
04030263FC731AE3
406282B300400293
005585B300550533
0032929340560633
0283839300000397
00038067405383B3
FE550EA3FFD58283
FE550F23FFE58283
FE550FA3FFF58283
02069863FC067693
FFC67693FA0600E3
00B68733F6068EE3
0005A28300367613
0055202300458593
FEE5E8E300450513
00B68733F5DFF06F
0005A28303F67613
0085A3830045A303
0105AE8300C5AE03
0185A8030145AF03
0055202301C5A883
0075242300652223
01D5282301C52623
01052C2301E52A23
0205A28301152E23
0285A3830245A303
0305AE8302C5AE03
0385A8030345AF03
0405859303C5A883
0265222302552023
03C5262302752423
03E52A2303D52823
03152E2303052C23
F6E5ECE304050513
00000000F41FF06F
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0200029300050F93
00060A6302567063
00B5002300A60733
FEE56CE300150513
00008067000F8513
0203006300357313
406282B300400293
4056063300550733
0015051300B50023
0FF5F593FEE51CE3
0055E5B300859293
0055E5B301059293
00367613FFC67693
03F6F29300A68733
FC05051300028E63
0000039700550533
405383B305038393
00B5202300038067
00B5242300B52223
00B5282300B52623
00B52C2300B52A23
02B5202300B52E23
02B5242302B52223
02B5282302B52623
02B52C2302B52A23
0405051302B52E23
F39FF06FFAE56EE3
0000000000000000
0000000000000000
0000000000000000
0000000000000000
0000000000000000
FF01011300000000
0121202300812423
1707879300000797
1684041300000417
0091222300112623
0287806340878933
0000049340295913
0014849300042783
000780E700440413
00000793FF24E8E3
0000009700078663
00000797000000E7
0000041712478793
4087893311C40413
00878E6340295913
0004278300000493
0044041300148493
FF24E8E3000780E7
0081240300C12083
0001290300412483
0000806701010113
00812423FF010113
0000079300112623
0007886300050413
0000009700000593
014000EF000000E7
088000EF00040513
0000806700050213
00812423FF010113
0987879300000797
0904041300000417
0091222340F40433
4024549300112623
FFC4041302048063
0004278300F40433
FFC40413FFF48493
FE0498E3000780E7
00078E6300000793
00C1208300812403
0101011300412483
0000006700000317
0081240300C12083
0101011300412483
FFFFF79700008067
00078C6354C78793
00100593FF010113
D34FF0EF00112623
0000006F0000006F
0000000000000000
0000000000000000
0000000400000000
0000000000000000
